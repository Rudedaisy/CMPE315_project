--
-- Entity: assign_0
-- Architecture : structural
-- Author: ehanson1
-- Created On: 10/28/2018
--
library STD;
library IEEE;
use IEEE.std_logic_1164.all;

entity assign_0 is

	port (
		output   : out std_logic);
end assign_0;

architecture structural of assign_0 is

begin

	output <= '0';

end structural;
